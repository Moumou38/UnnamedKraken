    ����          Assembly-CSharp   
PlayerData   	SceneNameCheckPointID	m_maxLifem_maxLightEnergym_maxJumpEnergym_coins           ReefBarrier                   